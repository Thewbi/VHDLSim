signal sinus_u     : unsigned(3 downto 0);