--Seconds + Minutes
--Seconds * 60
Seconds + Minutes * 60;