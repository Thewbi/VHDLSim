if rising_edge(clk) then
	q <= d;
end if;
