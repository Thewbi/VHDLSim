signal Counter : integer range 0 to 1;