--port map (a, b, c);
port map (d0, int_clk, q0);