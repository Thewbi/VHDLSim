use work.int_types.all;
