Y <= A OR B;