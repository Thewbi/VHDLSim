rising_edge(clk, a, b, c)