signal A : std_logic;