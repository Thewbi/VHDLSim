-- start symbol: alias_declaration

alias OpCode_s : bit_vector(7 downto 0) is Bus_s(31 downto 24);