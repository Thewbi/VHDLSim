if (bus_req_i.stb = '1') then
    rdata <= 1;
end if;