function Bitwise_AND (
    Seconds : integer := 0;
    a_vector : in std_logic_vector(3 downto 0);
    b_vector : out std_logic_vector(4 downto 1)
) return std_logic;

-- function Bitwise_AND (
--     Seconds : integer := 0;
--     a_vector : in std_logic_vector(3 downto 0);
--     b_vector : out std_logic_vector(4 downto 1)
-- );