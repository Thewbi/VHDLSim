-- start-symbol: if_statement

if OpCode_s = "10101011" then
    if Source_s = "1100" then
        Data16_s <= X"F904";
    end if;
end if;