type apples is range 0 to 100;
type oranges is range 0 to 100;

type day_of_month is range 0 to 31;
type year is range 0 to 2100;
