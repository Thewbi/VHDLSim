wait for 20 ns;