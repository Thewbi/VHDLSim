range 0 to CounterVal(Minutes => 1)