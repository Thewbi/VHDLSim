immediate <= replicate_f(exe_engine.ir(31), 21)