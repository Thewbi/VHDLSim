type t_FROM_FIFO is record
    wr_full  : std_logic;
    rd_empty : std_logic;
end record t_FROM_FIFO;