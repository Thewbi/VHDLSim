if rising_edge(clk, a, b, c) then
	q <= d;
end if;
