CounterVal(Minutes => 1) + 1