PACKAGE eight_bit_int IS 
    SUBTYPE BYTE IS INTEGER RANGE -128 TO 127; -- User-defined type
END eight_bit_int;