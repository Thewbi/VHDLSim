type resistance is range 0 to 1E9
units
    ohm;
end units resistance;
