signal rden  : std_ulogic;