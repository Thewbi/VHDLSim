read_ptr <= read_ptr + 1;