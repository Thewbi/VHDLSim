rden <= bus_req_i.stb and (not bus_req_i.rw);