entity flip.flap.flup.d_ff(basic)