--Seconds + Minutes
--Seconds * 60
--Seconds + Minutes * 60;
TotalSeconds * ClockFrequencyHz - 1;