--signal A : std_logic;

-- CounterVal() is a function
signal Counter : integer range 0 to CounterVal(Minutes => 1) + 1;