type alu_function is
 (disable, pass, add, subtract, multiply, divide);

type octal_digit is ('0', '1', '2', '3', '4', '5', '6', '7');
