-- start symbol: waveform_element

x"AB_CD_0955" after 10 ns;