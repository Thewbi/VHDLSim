Library IEEE;
use IEEE.std_logic_1164.all;

architecture orLogic of OR_gate is
begin
    Y <= A OR B;
end orLogic;