component OR_gate
    port (A : in std_logic;
          B : in std_logic;
          Y : out std_logic);
end component;