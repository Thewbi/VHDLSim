variable index : integer := 0;
variable sum, average, largest : real;
variable start, finish : time := 0 ns;
variable start : time := 0 ns; 
variable finish : time := 0 ns;
