bit0 : entity flip.flap.flup.d_ff(basic)
        port map (d0, int_clk, q0);